library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all

library work;

package global_package is
    type t_array_slv is array(natural range <>) of std_logic_vector;
end global_package;
